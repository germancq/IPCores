/**
 * @ Author: German Cano Quiveu, germancq
 * @ Create Time: 2020-01-19 13:34:50
 * @ Modified by: Your name
 * @ Modified time: 2020-02-19 11:37:46
 * @ Description:
 */

 package configuration;
    loclparam CLK_INTERNAL_DIVIDER = 17
    loclparam N_BLOCK_SIZE = 32,
    loclparam SCLK_SPEED_SIZE = 5,
    loclparam CMD18_SIZE = 1,
    loclparam START_BLOCK = 32'h0x00100000

endpackage