/**
 * @ Author: German Cano Quiveu, germancq
 * @ Create Time: 2020-01-19 13:34:50
 * @ Modified by: germancq
 * @ Modified time: 2020-01-19 13:44:17
 * @ Description:
 */

 package configuration;
    loclparam CLK_INTERNAL_DIVIDER = 17
    loclparam SIZE_OUTPUT_UUT_1 = 8,
    loclparam SIZE_OUTPUT_UUT_2 = 8,
    loclparam SIZE_INPUT_UUT_1 = 32,
    loclparam START_BLOCK = 32'h0x00100000

endpackage